module singlecycle_tb;

logic [
